// reloj_soc_tb.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module reloj_soc_tb (
	);

	wire         reloj_soc_inst_clk_bfm_clk_clk;            // reloj_soc_inst_clk_bfm:clk -> [reloj_soc_inst:clk_clk, reloj_soc_inst_reset_bfm:clk]
	wire   [7:0] reloj_soc_inst_buttons_bfm_conduit_export; // reloj_soc_inst_buttons_bfm:sig_export -> reloj_soc_inst:buttons_export
	wire  [31:0] reloj_soc_inst_leds_export;                // reloj_soc_inst:leds_export -> reloj_soc_inst_leds_bfm:sig_export
	wire         reloj_soc_inst_reset_bfm_reset_reset;      // reloj_soc_inst_reset_bfm:reset -> reloj_soc_inst:reset_reset_n

	reloj_soc reloj_soc_inst (
		.buttons_export (reloj_soc_inst_buttons_bfm_conduit_export), // buttons.export
		.clk_clk        (reloj_soc_inst_clk_bfm_clk_clk),            //     clk.clk
		.leds_export    (reloj_soc_inst_leds_export),                //    leds.export
		.reset_reset_n  (reloj_soc_inst_reset_bfm_reset_reset)       //   reset.reset_n
	);

	altera_conduit_bfm reloj_soc_inst_buttons_bfm (
		.sig_export (reloj_soc_inst_buttons_bfm_conduit_export)  // conduit.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) reloj_soc_inst_clk_bfm (
		.clk (reloj_soc_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm_0002 reloj_soc_inst_leds_bfm (
		.sig_export (reloj_soc_inst_leds_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) reloj_soc_inst_reset_bfm (
		.reset (reloj_soc_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (reloj_soc_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
